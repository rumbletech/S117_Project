library verilog;
use verilog.vl_types.all;
entity SPI_TB is
end SPI_TB;
